module main

fn test_collatz() {
	assert collatz(13) == 9
}
